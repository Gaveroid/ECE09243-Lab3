module Decoder(select, enable, x);

	input [4:0] select;
	input enable;
	
	output reg [31:0] x;
	
	always @(select)
	begin
		if (enable==1)
			case (select)
				5'd0: x <= 32'b00000000000000000000000000000001;
				5'd1: x <= 32'b00000000000000000000000000000010;
				5'd2: x <= 32'b00000000000000000000000000000100;
				5'd3: x <= 32'b00000000000000000000000000001000;
				5'd4: x <= 32'b00000000000000000000000000010000;
				5'd5: x <= 32'b00000000000000000000000000100000;
				5'd6: x <= 32'b00000000000000000000000001000000;
				5'd7: x <= 32'b00000000000000000000000010000000;
				5'd8: x <= 32'b00000000000000000000000100000000;
				5'd9: x <= 32'b00000000000000000000001000000000;
				5'd10: x <= 32'b00000000000000000000010000000000;
				5'd11: x <= 32'b00000000000000000000100000000000;
				5'd12: x <= 32'b00000000000000000001000000000000;
				5'd13: x <= 32'b00000000000000000010000000000000;
				5'd14: x <= 32'b00000000000000000100000000000000;
				5'd15: x <= 32'b00000000000000001000000000000000;
				5'd16: x <= 32'b00000000000000010000000000000000;
				5'd17: x <= 32'b00000000000000100000000000000000;
				5'd18: x <= 32'b00000000000001000000000000000000;
				5'd19: x <= 32'b00000000000010000000000000000000;
				5'd20: x <= 32'b00000000000100000000000000000000;
				5'd21: x <= 32'b00000000001000000000000000000000;
				5'd22: x <= 32'b00000000010000000000000000000000;
				5'd23: x <= 32'b00000000100000000000000000000000;
				5'd24: x <= 32'b00000001000000000000000000000000;
				5'd25: x <= 32'b00000010000000000000000000000000;
				5'd26: x <= 32'b00000100000000000000000000000000;
				5'd27: x <= 32'b00001000000000000000000000000000;
				5'd28: x <= 32'b00010000000000000000000000000000;
				5'd29: x <= 32'b00100000000000000000000000000000;
				5'd30: x <= 32'b01000000000000000000000000000000;
				5'd31: x <= 32'b10000000000000000000000000000000;
			endcase
			else if (enable==0) x <= 32'b00000000000000000000000000000000;
	end
	
endmodule
